`timescale 1ns / 1ps

module Cactus(
    input wire [31:0] clkdiv,
    input wire RESET,
    input wire START,
    input wire [8:0] row_addr,
    input wire [9:0] col_addr,
    input wire game_status,
    input wire fresh,
    input wire [3:0] speed,
    output reg px
    );

    reg [59:0] pattern [57:0];
    reg [9:0] position;


    always @(negedge fresh) begin
        if (game_status) begin
            position<=(position+speed)%(10'd640+10'd60);
        end else begin
            if (RESET || START) begin
                position <=10'b0;
            end
        end
    end

    always @(posedge clkdiv[0]) begin
        //TEST
        // if (game_status) begin
            if (row_addr>=10'd344 && row_addr<10'd402) begin
                if (col_addr>=(10'd640 > position ? 10'd640 - position : 10'd0) && col_addr<10'd700 - position) begin
                    px <= pattern[row_addr - 16'd344][col_addr + position - 16'd640];
                end else begin
                    px <= 1'b0;
                end
            end else begin
                px <= 1'b0;
            end
        // end
    end


    always @(posedge RESET) begin
        //row 58
        //col 60
        pattern[0]<=60'b0000000000_0000000000_0000000111_1110000000_0000000000_0000000000;
        pattern[1]<=60'b0000000000_0000000000_0000001111_1111000000_0000000000_0000000000;
        pattern[2]<=60'b0000000000_0000000000_0000011111_1111100000_0000000000_0000000000;
        pattern[3]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[4]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[5]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[6]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[7]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[8]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[9]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[10]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[11]<=60'b0000000000_0000011000_0000111111_1111110000_0000000000_0000000000;
        pattern[12]<=60'b0000000000_0000111100_0000111111_1111110000_0000000000_0000000000;
        pattern[13]<=60'b0000000000_0001111110_0000111111_1111110000_0000000000_0000000000;
        pattern[14]<=60'b0000000000_0011111111_0000111111_1111110000_0011000000_0000000000;
        pattern[15]<=60'b0000000000_0011111111_0000111111_1111110000_0111100000_0000000000;
        pattern[16]<=60'b0000000000_0011111111_0000111111_1111110000_1111110000_0000000000;
        pattern[17]<=60'b0000000000_0011111111_0000111111_1111110000_1111110000_0000000000;
        pattern[18]<=60'b0000000000_0011111111_0000111111_1111110000_1111110000_0000000000;
        pattern[19]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        pattern[20]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        pattern[21]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        pattern[22]<=60'b0000000000_0011111111_1111111111_1111110000_1111110000_0000000000;
        pattern[23]<=60'b0000000000_0011111111_1111111111_1111111111_1111110000_0000000000;
        pattern[24]<=60'b0000000000_0000111111_1111111111_1111111111_1111110000_0000000000;
        pattern[25]<=60'b0000000000_0000001111_1111111111_1111111111_1111110000_0000000000;
        pattern[26]<=60'b0000000000_0000000011_1111111111_1111111111_1111000000_0000000000;
        pattern[27]<=60'b0000000000_0000000000_1111111111_1111111111_1100000000_0000000000;
        pattern[28]<=60'b0000000000_0000000000_0000111111_1111111111_0000000000_0000000000;
        pattern[29]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[30]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[31]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[32]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[33]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[34]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[35]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[36]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[37]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[38]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[39]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[40]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[41]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[42]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[43]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[44]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[45]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[46]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[47]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[48]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[49]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[50]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[51]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[52]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[53]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[54]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[55]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[56]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
        pattern[57]<=60'b0000000000_0000000000_0000111111_1111110000_0000000000_0000000000;
    end
    

endmodule
