`timescale 1ns / 1ps

module Cactus(
    input wire [31:0] clkdiv,
    input wire [8:0] row_addr,
    input wire [9:0] col_addr,
    output reg [9:0] ground_position,
    input wire game_status,
    input wire fresh,
    input wire [3:0] speed,
    output reg px
    );
    
    
    

endmodule
