`timescale 1ns / 1ps

module Jump (
    input wire fresh,
    input wire [31:0] clkdiv,
    input wire button_jump,
    input wire RESET,
    input wire START,
    input wire [8:0] row_addr,
    input wire [9:0] col_addr,
    output reg px,
    input wire game_status
    );
    
    reg [11:0] jump_time;
    wire [11:0] height;
    reg [0:82] body_run [0:73];
    reg [0:82] body_stop [0:73];
    reg [0:82] feet_stop [0:13];
    reg [0:82] feet_run_a [0:13];
    reg [0:82] feet_run_b [0:13];
    reg jumping;

    reg [3:0] counter;

    //height is only associated with the value of jump_time
    assign height = (jump_time*12'd40 - jump_time*jump_time) / 2'd2;

    //for every frame
    always @(negedge fresh) begin //negedge guarantees the operation are done in the blanking period
        //add counter
        counter<=counter+1;
        //jump operation
        if (game_status) begin
            if (button_jump && jumping==1'b0) begin
               jumping<=1'b1;//begin to jump
            end
            if (jumping) begin
                if (jump_time>=12'd40) begin//reset jump operation
                    jump_time<=12'b0;
                    jumping<=1'b0;
                end else begin
                    jump_time<=jump_time+1'b1;//add jump_time
                end
            end
        end else begin //if pausing
            if (RESET || START) begin
                jump_time<=12'b0;
                jumping<=1'b0;
                counter<=4'b0;
            end
            //if neither RESET nor START, do nothing to keep the current position of the dinosaur
        end
        
    end

    always @(posedge clkdiv[0]) begin
        //caculate the value of px based on row_addr and col_addr
        //body part
        if (row_addr >= 10'd402 - height - 10'd88 && row_addr < 10'd402 - height -10'd14 && col_addr>=10'd80 && col_addr<10'd162) begin
            if (game_status) begin //if running
                px <= body_run[row_addr+height-10'd314][col_addr-12'd80];
            end else begin //if it stops
                px <= body_stop[row_addr+height-10'd314][col_addr-12'd80];
            end
            
        end else begin
            px <= 1'b0;
        end

        //feet part
        if (row_addr >= 10'd402 - height - 10'd14 && row_addr < 10'd402 - height && col_addr>=10'd80 && col_addr<10'd162) begin
            if (game_status && height==0) begin
                //moving feet
                if (counter[3]) begin
                    px<=feet_run_a[row_addr+height-10'd388][col_addr-12'd80];
                end else begin
                    px<=feet_run_b[row_addr+height-10'd388][col_addr-12'd80];
                end
            end else begin
                //stopped feet
                px<=feet_stop[row_addr+height-10'd388][col_addr-12'd80];
            end

        end

    end

    always @(posedge RESET) begin
        //use ram to store the pattern of dinosaur (row 88, col 82)
        body_run[0]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_run[1]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_run[2]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_run[3]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_run[4]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[5]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[6]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[7]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[8]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1100011111_1111111111_1111111111_11;
        body_run[9]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1100011111_1111111111_1111111111_11;
        body_run[10]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1100011111_1111111111_1111111111_11;
        body_run[11]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[12]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[13]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[14]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[15]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[16]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[17]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[18]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[19]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[20]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[21]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[22]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_run[23]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1110000000_0000000000_00;
        body_run[24]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1110000000_0000000000_00;
        body_run[25]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1110000000_0000000000_00;
        body_run[26]<=82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
        body_run[27]<=82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
        body_run[28]<=82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[29]<=82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[30]<=82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[31]<=82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[32]<=82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[33]<=82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[34]<=82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[35]<=82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[36]<=82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[37]<=82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[38]<=82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_run[39]<=82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_run[40]<=82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_run[41]<=82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_run[42]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_run[43]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_run[44]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_run[45]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_run[46]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[47]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[48]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[49]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[50]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[51]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[52]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[53]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[54]<=82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[55]<=82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[56]<=82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[57]<=82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[58]<=82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[59]<=82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[60]<=82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[61]<=82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_run[62]<=82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
        body_run[63]<=82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
        body_run[64]<=82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
        body_run[65]<=82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
        body_run[66]<=82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
        body_run[67]<=82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
        body_run[68]<=82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
        body_run[69]<=82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
        body_run[70]<=82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
        body_run[71]<=82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
        body_run[72]<=82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
        body_run[73]<=82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;


        feet_stop[0]<=82'b0000000000_0000000000_1111111111_1100001111_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[1]<=82'b0000000000_0000000000_1111111111_1100001111_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[2]<=82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[3]<=82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[4]<=82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[5]<=82'b0000000000_0000000000_1111110000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[6]<=82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[7]<=82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[8]<=82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[9]<=82'b0000000000_0000000000_1111000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_stop[10]<=82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
        feet_stop[11]<=82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
        feet_stop[12]<=82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;
        feet_stop[13]<=82'b0000000000_0000000000_1111111100_0000000000_1111111100_0000000000_0000000000_0000000000_00;


        feet_run_a[0]<=82'b0000000000_0000000000_1111111100_0000001111_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[1]<=82'b0000000000_0000000000_1111111100_0000001111_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[2]<=82'b0000000000_0000000000_1111111100_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[3]<=82'b0000000000_0000000000_0011111111_1111000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[4]<=82'b0000000000_0000000000_0011111111_1111000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[5]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[6]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[7]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[8]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[9]<=82'b0000000000_0000000000_0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_a[10]<=82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
        feet_run_a[11]<=82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
        feet_run_a[12]<=82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;
        feet_run_a[13]<=82'b0000000000_0000000000_0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_00;


        feet_run_b[0]<=82'b0000000000_0000000000_1111111111_1100000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_b[1]<=82'b0000000000_0000000000_1111111111_1100000000_1111000000_0000000000_0000000000_0000000000_00;
        feet_run_b[2]<=82'b0000000000_0000000000_1111111100_0000000000_1111111111_0000000000_0000000000_0000000000_00;
        feet_run_b[3]<=82'b0000000000_0000000000_1111111100_0000000000_1111111111_0000000000_0000000000_0000000000_00;
        feet_run_b[4]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_run_b[5]<=82'b0000000000_0000000000_1111110000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_run_b[6]<=82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_run_b[7]<=82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_run_b[8]<=82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_run_b[9]<=82'b0000000000_0000000000_1111000000_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_run_b[10]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_run_b[11]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_run_b[12]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;
        feet_run_b[13]<=82'b0000000000_0000000000_1111111100_0000000000_0000000000_0000000000_0000000000_0000000000_00;



        body_stop[0]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_stop[1]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_stop[2]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_stop[3]<=82'b0000000000_0000000000_0000000000_0000000000_0000000011_1111111111_1111111111_1111111100_00;
        body_stop[4]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[5]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[6]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
        body_stop[7]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
        body_stop[8]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0011001111_1111111111_1111111111_11;
        body_stop[9]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0011001111_1111111111_1111111111_11;
        body_stop[10]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
        body_stop[11]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_0000001111_1111111111_1111111111_11;
        body_stop[12]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[13]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[14]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[15]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[16]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[17]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[18]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[19]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[20]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[21]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[22]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[23]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111111_11;
        body_stop[24]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111100_00;
        body_stop[25]<=82'b0000000000_0000000000_0000000000_0000000000_0000111111_1111111111_1111111111_1111111100_00;
        body_stop[26]<=82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
        body_stop[27]<=82'b1111000000_0000000000_0000000000_0000000000_1111111111_1111111111_1111111111_1111111100_00;
        body_stop[28]<=82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[29]<=82'b1111000000_0000000000_0000000000_0000001111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[30]<=82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[31]<=82'b1111000000_0000000000_0000000000_0000111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[32]<=82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[33]<=82'b1111110000_0000000000_0000000000_0011111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[34]<=82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[35]<=82'b1111111100_0000000000_0000000000_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[36]<=82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[37]<=82'b1111111111_0000000000_0000001111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[38]<=82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_stop[39]<=82'b1111111111_1100000000_0000111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_stop[40]<=82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_stop[41]<=82'b1111111111_1111000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_00;
        body_stop[42]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_stop[43]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_stop[44]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_stop[45]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_1111000000_0000000000_00;
        body_stop[46]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[47]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[48]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[49]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[50]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[51]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[52]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[53]<=82'b1111111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[54]<=82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[55]<=82'b0011111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[56]<=82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[57]<=82'b0000111111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[58]<=82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[59]<=82'b0000001111_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[60]<=82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[61]<=82'b0000000011_1111111111_1111111111_1111111111_1111111111_1111110000_0000000000_0000000000_00;
        body_stop[62]<=82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
        body_stop[63]<=82'b0000000000_1111111111_1111111111_1111111111_1111111111_1111000000_0000000000_0000000000_00;
        body_stop[64]<=82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
        body_stop[65]<=82'b0000000000_0011111111_1111111111_1111111111_1111111111_1100000000_0000000000_0000000000_00;
        body_stop[66]<=82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
        body_stop[67]<=82'b0000000000_0000111111_1111111111_1111111111_1111111111_0000000000_0000000000_0000000000_00;
        body_stop[68]<=82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
        body_stop[69]<=82'b0000000000_0000001111_1111111111_1111111111_1111111100_0000000000_0000000000_0000000000_00;
        body_stop[70]<=82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
        body_stop[71]<=82'b0000000000_0000000011_1111111111_1111111111_1111110000_0000000000_0000000000_0000000000_00;
        body_stop[72]<=82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
        body_stop[73]<=82'b0000000000_0000000000_1111111111_1111111111_1111000000_0000000000_0000000000_0000000000_00;
      end
    
 
    
endmodule
